* # FILE NAME: /HOME/ECEGRID/A/559MG3/CADENCE/SIMULATION/CMOS_NAND_180NM/       
* HSPICES/EXTRACTED/NETLIST/CMOS_NAND_180NM.C.RAW
* NETLIST OUTPUT FOR HSPICES.
* GENERATED ON OCT 31 15:04:53 2014
   
* FILE NAME: HW1_CMOS_NAND_180NM_EXTRACTED.S.
* SUBCIRCUIT FOR CELL: CMOS_NAND_180NM.
* GENERATED FOR: HSPICES.
* GENERATED ON OCT 31 15:04:53 2014.
   
M2 VDD! B OUT VDD!  TSMC18DP  L=180.000000682412E-9 W=810.000017281709E-9 
+AD=364.499988352029E-15 AS=218.700003853239E-15 PD=1.70999999227206E-6 
+PS=539.999973625527E-9 M=1 
M3 OUT A VDD! VDD!  TSMC18DP  L=180.000000682412E-9 W=810.000017281709E-9 
+AD=218.700003853239E-15 AS=364.499988352029E-15 PD=539.999973625527E-9 
+PS=1.70999999227206E-6 M=1 
M4 OUT B 1 0  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=251.100003420199E-15 AS=72.8999990256586E-15 PD=2.06999993679347E-6 
+PS=539.999973625527E-9 M=1 
M5 1 A 0 0  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=72.8999990256586E-15 AS=226.799996968716E-15 PD=539.999973625527E-9 
+PS=1.89000002137618E-6 M=1 
   
   
   
   
   
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc18dP" PMOS 
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc18dN" NMOS 
   
   
* INCLUDE FILES
   
   
 
   
* END OF NETLIST
.TEMP    25.0000    
*.OP
*.save
*.OPTION  INGOLD=2 ARTIST=2 PSF=2
*+        PROBE=0
vvdd! vdd! 0 DC=2.5v
.END
