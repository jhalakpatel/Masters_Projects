* # FILE NAME: /HOME/ECEGRID/A/559MG3/CADENCE/SIMULATION/INVERTERTEST/          
* HSPICES/SCHEMATIC/NETLIST/INVERTERTEST.C.RAW
* NETLIST OUTPUT FOR HSPICES.
* GENERATED ON OCT 18 21:13:12 2014
   
* GLOBAL NET DEFINITIONS
.GLOBAL VDD! 
* FILE NAME: JHALAK_LIB_INVERTERTEST_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: INVERTERTEST.
* GENERATED FOR: HSPICES.
* GENERATED ON OCT 18 21:13:12 2014.
.SUBCKT InverterTest IN_0 IN_1 OUT_0 OUT_1  
XI9 IN_0 INTERNAL_0 INVERTERP_1 
XI10 IN_1 NET21 INVERTERP_1 
XI14 NET21 INTERNAL_1 INVERTERP_1 
XI12 INTERNAL_1 OUT_1 INVERTERP_1 
XI13 INTERNAL_0 OUT_0 INVERTERP_1 
C1 OUT_0 0  10E-15 M=1.0 
C0 OUT_1 0  10E-15 M=1.0 
.ENDS

* FILE NAME: JHALAK_LIB_INVERTERP_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: INVERTERP.
* GENERATED FOR: HSPICES.
* GENERATED ON OCT 18 21:13:12 2014.
   
* TERMINAL MAPPING: IN = IN
*                   OUT = OUT
.SUBCKT INVERTERP_1 IN OUT 
MP0 OUT IN VDD! VDD!  TSMC25P  L=(2.4E-07) W=(6E-07) AD=+4.50000000E-13 
+AS=+4.50000000E-13 PD=+2.70000000E-06 PS=+2.70000000E-06 M=1 
MN0 OUT IN 0 0  TSMC25N  L=(2.4E-07) W=(3E-07) AD=+2.25000000E-13 
+AS=+2.25000000E-13 PD=+2.10000000E-06 PS=+2.10000000E-06 M=1 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS INVERTERP_1 
   
   
   
   
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc25N" NMOS 
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc25P" PMOS 
   
* INCLUDE FILES
   
   
   
   
   
   
* END OF NETLIST
.TRAN  1.00000E-09 3.00000E-08 START=  0.0000    
.TEMP    25.0000    
.OP
.save
.OPTION  INGOLD=2 ARTIST=2 PSF=2
+        PROBE=0
vin_1 in_1 0 pulse 0.0 2.5 1n 1n 1n 10n 20n
vin_0 in_0 0 pulse 0.0 2.5 1n 1n 1n 10n 20n
vvdd! VDD! 0 DC=2.5v
.END
