* # FILE NAME: /HOME/ECEGRID/A/559MG3/CADENCE/SIMULATION/CMOS_NOR_180NM/        
* HSPICES/SCHEMATIC/NETLIST/CMOS_NOR_180NM.C.RAW
* NETLIST OUTPUT FOR HSPICES.
* GENERATED ON OCT 31 14:54:14 2014
   
* GLOBAL NET DEFINITIONS
.GLOBAL VDD! 
* FILE NAME: HW1_CMOS_NOR_180NM_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: CMOS_NOR_180NM.
* GENERATED FOR: HSPICES.
* GENERATED ON OCT 31 14:54:14 2014.
   
MP0 OUT A NET11 VDD!  TSMC18DP  L=180E-9 W=810E-9 AD=364.5E-15 AS=364.5E-15 
+PD=2.52E-6 PS=2.52E-6 M=1 
MP1 NET11 B VDD! VDD!  TSMC18DP  L=180E-9 W=810E-9 AD=364.5E-15 AS=364.5E-15 
+PD=2.52E-6 PS=2.52E-6 M=1 
MN0 OUT A 0 0  TSMC18DN  L=180E-9 W=270E-9 AD=121.5E-15 AS=121.5E-15 
+PD=1.44E-6 PS=1.44E-6 M=1 
MN1 OUT B 0 0  TSMC18DN  L=180E-9 W=270E-9 AD=121.5E-15 AS=121.5E-15 
+PD=1.44E-6 PS=1.44E-6 M=1 
   
   
   
   
   
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc18dP" PMOS 
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc18dN" NMOS 
   
   
* INCLUDE FILES
   
   
   
   
   
   
* END OF NETLIST
.TEMP    25.0000    
*.OP
*.save
*.OPTION  INGOLD=2 ARTIST=2 PSF=2
*+        PROBE=0
vvdd! vdd! 0 DC=2.5v
.END
